`timescale 1ps/1ps
`define DATA_WIDTH 4
`define N 3

module balanced_adder_tb ();

	// note this only runs for 50 cycles with the below settings
	// alter TB_TIMEOUT to run longer
	localparam TB_TIMEOUT    = 100000;
	localparam TB_CLK_PERIOD = 2000;
	localparam TB_RST_PERIOD = 4000;

	initial  #(TB_TIMEOUT) $finish();

	// clock
	reg tb_clk = 1'b0;
	always #(TB_CLK_PERIOD/2) tb_clk = ~tb_clk;
//reg[10:0] k;

	// DUT
	wire [`DATA_WIDTH*`N-1 : 0] outp;
	wire [`DATA_WIDTH*(2**`N) - 1 : 0] inps;


	balanced_adder_test #(
		.data_width(`DATA_WIDTH),
                .N(`N)
	) my_adder (
		.clk(tb_clk),
		.outp(outp),
		.outp_inps(inps)
		);
	// display inputs and output on each clock cycle
	always @(posedge tb_clk) begin
		$display("inps = ", inps, " => outp = ", outp);
     //     for (k = 1; k <= 2**(N-1); k = k + 1) begin
		//$display("inps = ", inps[k*`DATA_WIDTH-1:(k-1)*`DATA_WIDTH], " => outp = ", outp);

      //    end     

	end

endmodule
